//------------------------------------------------
// mipsmem.v
// David_Harris@hmc.edu 23 October 2005
// External memories used by MIPS processors
//------------------------------------------------


module dmem(input         clk, we,
            input  [31:0] a, wd,
            output [31:0] rd);

  reg  [31:0] RAM[63:0];

  always @(posedge clk)
    if (we)
      RAM[a[31:2]] <= wd;
  assign rd = RAM[a[31:2]]; // word aligned
endmodule


